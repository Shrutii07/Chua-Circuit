*Chua OPAMP

.include LF356.MOD
V1 2 0 dc 9
V2 5 0 dc -9

L 1 0 18m
C1 1 0 100n
C2 9 0 10n
R 1 9 1.6K

XU1 9 4 2 5 6 LF356/NS
XU2 9 7 2 5 8 LF356/NS
R1 8 9 22K
R2 8 7 22K
R3 7 0 3.3K
R4 6 9 220
R5 6 4 220
R6 4 0 2.2K


.tran 1u 10m
.control

SET COLOR0 = white
SET COLOR1 = black
SET COLOR2= red
SET COLOR3= blue
SET COLOR4 = brown
Set XbrushWidth = 2

run
.options savecurrents
*plot -(@R4[i]+@R1[i]) vs V(9)
plot v(1) vs v(9)
*plot v(1) v(9)
*plot V(1) V(9)
*linearize
*fft V(1) V(9)
*plot V(1) V(9) xlimit 0 10kHz
.endc
.end
